`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name:    instr_mem 
//////////////////////////////////////////////////////////////////////////////////
module instr_mem     
 (  
      input     [31:0]     pc,  
      output wire     [31:0]          instruction  
 );  
      wire [4 : 0] rom_addr;
      //assign rom_addr = pc[4 : 1];  
      assign rom_addr = pc[4 : 0];
      reg [31:0] rom[31:0];  
      initial  
      begin  
                rom[0] = 32'b00000000000000000000000000000000;
                rom[1] = 32'b00000000001000100001100000000000; //add
			 rom[2] = 32'b00000000100001010011000000000000; //ADD
                rom[3] = 32'b00011000111001110000000000000111; // branch equal 
                //rom[3] = 32'b00000000111010000100100000000000; //add
                rom[4] = 32'b00000001010010110110000000000000; //add
			 rom[5] = 32'b00000001101011100111100000000000; //ADD
                rom[6] = 32'b00000010000100011001000000000000; //add
                //rom[3] = 32'b00000000111001100000100000000001; //SUB					 
                //rom[4] = 32'b00011100111001100000000000000111; //ADI
                //rom[5] = 32'b00000000111001100000000000000010; //AND
                rom[7] = 32'b00000010011101001010100000000000; //add
			 rom[8] = 32'b00000010110101111100000000000000; //ADD
                rom[9] = 32'b00000011001110101101100000000000; //add
                rom[10] = 32'b00000011100111011111000000000000; //add
			 rom[11] = 32'b00000000001000110010000000000000; //ADD
                rom[12] = 32'b00000000111010000100100000000000; //add					 
                rom[13] = 32'b00000001010010110110000000000000;  //add 
                rom[14] = 32'b00000001100011100111100000000000;  //add hazard
                rom[15] = 32'b00000010000100011001000000000000; //add
                rom[16] = 32'b00001000000000000000000000000111; // jump 
                rom[17]= 32'b00011000111001100000000000000100; //SLT
                rom[18]= 32'b00000000111000010011000000001000; //jr
                rom[19]= 32'b00000000111000010011000000001000;  
                rom[20]= 32'b00010000010000110000000000000000;  //ld 
                //$finish;
      end  
      assign instruction = (pc[31:0] < 32 )? rom[rom_addr[4:0]]: 32'd0; 
       
 endmodule   
