`timescale 1ns / 1ps
package spi_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "../uvm/spi_sequence_item.sv"
`include "../uvm/spi_sequence.sv"
`include "../uvm/spi_driver.sv"
`include "../uvm/spi_interface.sv"
`include "../uvm/spi_monitor.sv"
`include "../uvm/spi_agent.sv"
`include "../uvm/spi_scorecard.sv"
`include "../uvm/spi_environment.sv"
`include "../uvm/spi_test.sv"

    
endpackage